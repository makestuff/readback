lx9r1.vhdl